grammar edu:umn:cs:melt:exts:ableC:regexInADT:mda_test;

import edu:umn:cs:melt:exts:ableC:algDataTypes:artifact;

copper_mda testPatternRegex(extendedParser) {
  edu:umn:cs:melt:exts:ableC:regexInADT;
}

